----------------------------------------------------------------------------------

-- Group 17
-- Senevirathne S.M.P.U.
-- 
-- Create Date: 04/16/2024 02:13:42 PM
-- Design Name: Carry_Look_Ahead_Adder_Subtractor
-- Module Name: Carry_Look_Ahead_Adder_Subtractor - Behavioral
-- Project Name: Nanoprocessor
-- Target Devices: Basys3 Board

----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Carry_Look_Ahead_Adder_Subtractor is
    Port ( A : in STD_LOGIC_VECTOR (3 downto 0); --Bus for the first binary number
           B : in STD_LOGIC_VECTOR (3 downto 0); --Bus for the second binary number
           Add_Sub : in STD_LOGIC; --Should we add B to A or should we subtract B from A? (1 for subtraction, 0 for addition)
           EN : in STD_LOGIC; --Enable input
           S : inout STD_LOGIC_VECTOR (3 downto 0); --Bus for the binary sum output
           Sign : inout STD_LOGIC; --Sign Bit: 1 for negative, 0 for positive
           Overflow : inout STD_LOGIC; --Overflow bit: Is there an overflow?
           --When the number is negative, is the number in range [-0,-8]: if yes, there is no overflow => Overflow =0; if no, there is an overflow => Overflow = 1
           --When the number is positive, is the number in range [+0, 7]: if yes, there is no overflow => Overflow =0; if no, there is an overflow => Overflow = 1
           Zero : inout STD_LOGIC); --Is the output zero(0000) even when Enable is 1?
end Carry_Look_Ahead_Adder_Subtractor;

architecture Behavioral of Carry_Look_Ahead_Adder_Subtractor is
component Full_Adder is
    Port ( A : in STD_LOGIC; --First input bit
           B : in STD_LOGIC; --Second input bit
           Carry_in : in STD_LOGIC; --Carry input bit
           Sum : out STD_LOGIC; --Sum output bit
           Carry_out : out STD_LOGIC; --Carry output bit
           P : out STD_LOGIC; --Propergate output bit
           G : out STD_LOGIC); --Generate output bit
end component;

component Carry_Look_Ahead is
    Port ( P : in STD_LOGIC_VECTOR (2 downto 0); --Propergate input bus
           G : in STD_LOGIC_VECTOR (2 downto 0); --Propergate output bus
           Carry_in : in STD_LOGIC; --Carry input bit
           Carry_out : out STD_LOGIC_VECTOR (3 downto 2)); --Carry output bus
end component;

--Signal the inputs and outputs of internal components
SIGNAL A0, B0, C1, P0, G0: std_logic; --FA0
SIGNAL A1, B1, P1, G1: std_logic; --FA1
SIGNAL A2, B2, C2, P2, G2: std_logic; --FA2
SIGNAL A3, B3, C3, C4: std_logic; --FA3

--An and Bn are n th bits of the binary numbers A and B inserted to the relevant(n th) Full Adder
--Cn is the carry bit generated by adding the n th bits of A and B
--Pn and Gn are propergation and generation bits of the relevant(n th) Full Adder
begin
    Full_Adder_0 : Full_Adder --mapping first full adder
        port map(A => A0,
        B => B0,
        Carry_in => Add_Sub, --C0
        Sum => S(0),
        Carry_out => C1,
        P => P0,
        G => G0
    );
    Full_Adder_1 :Full_Adder --mapping second full adder
        port map(A => A1,
        B => B1,
        Carry_in => C1,
        Sum => S(1),
        P => P1,
        G => G1
    );
    Full_Adder_2 :Full_Adder --mapping third full adder
        port map(A => A2,
        B => B2,
        Carry_in => C2,
        Sum => S(2),
        P => P2,
        G => G2
    );
    Full_Adder_3 :Full_Adder --mapping last full adder
        port map(A => A3,
        B => B3,
        Carry_in => C3,
        Sum => S(3),
        Carry_out => C4 
    );
    Carry_Look_Ahead_0 : Carry_Look_Ahead --mapping carry look ahead logic unit
        port map(P(0) => P0, P(1) => P1, P(2) => P2,
        G(0) => G0, G(1) => G1, G(2) => G2,
        Carry_in => Add_Sub, --C0
        Carry_out(2) => C2, Carry_out(3) => C3
    );

--Defining inputs of FA0 (A0, B0)
A0 <= (EN AND A(0)) XOR Add_Sub;
B0 <= B(0) AND EN;

--Defining inputs of FA1 (A1, B1)
A1 <= (EN AND A(1)) XOR Add_Sub;
B1 <= B(1) AND EN;

--Defining inputs of FA2 (A2, B2)
A2 <= (EN AND A(2)) XOR Add_Sub;
B2 <= B(2) AND EN;

--Defining inputs of FA3 (A3, B3)
A3 <= (EN AND A(3)) XOR Add_Sub;
B3 <= B(3) AND EN;

--Defining the zero flag
Zero <= EN AND NOT(S(0) OR S(1) OR S(2) OR S(3));

--carry output of the Carry Look Ahead Adder Subtractor
Sign <= (S(3) AND NOT(Overflow)) OR (NOT(A(3)) AND Overflow AND Add_Sub);

--Defining the overflow bit
Overflow <= C3 XOR (C4 );

end Behavioral;
